package afvip_pkg;
  import uvm_pkg::*;


	`include "uvm_macros.svh"
	`include "afvip_item.svh"
    `include "afvip_sequencer.svh"
	`include "afvip_driver.svh"
	`include "afvip_monitor.svh"
	`include "afvip_agent.svh"
	`include "afvip_sequence.svh"
	`include "afvip_coverage.svh"

endpackage : afvip_pkg;