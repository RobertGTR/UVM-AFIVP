package tb_pkg;
import uvm_pkg::*;
import afvip_pkg::*;
import interr_pkg::*;
import reset_pkg::*;

 `include "uvm_macros.svh"
 `include "my_scoreboard.svh"
 `include "afvip_env.svh"
 `include "afvip_test.svh"

endpackage:tb_pkg
 