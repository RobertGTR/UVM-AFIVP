package interr_pkg;
      import uvm_pkg::*;

   `include "uvm_macros.svh"
   `include "afvip_interrupt_item.svh"
   `include "afvip_interrupt_monitor.svh"
   `include "afvip_interrupt_agent.svh"

endpackage:interr_pkg
